interface mux_if; 
  logic [3:0] in0; 
  logic [3:0] in1; 
  logic [3:0] in2; 
  logic [3:0] in3; 
  logic [1:0] sel; 
  logic [3:0] out; 
endinterface
  